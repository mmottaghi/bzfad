
`timescale 1 ns/10 ps
module evRst_Latch_cell_5 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evRst_Latch_cell_4 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evRst_Latch_cell_3 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evRst_Latch_cell_2 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evRst_Latch_cell_1 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evRst_Latch_cell_0 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evCINV_30 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_29 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_28 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_27 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_26 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_25 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_24 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_23 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_22 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_21 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_20 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_19 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_18 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_17 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_16 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_15 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_14 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_13 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_12 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_11 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_10 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_9 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_8 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_7 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_6 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_5 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_4 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_3 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_2 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_1 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evCINV_0 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_30 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_29 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_28 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_27 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_26 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_25 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_24 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_23 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_22 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_21 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_20 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_19 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_18 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_17 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_16 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_15 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_14 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_13 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_12 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_11 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_10 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_9 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_8 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_7 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_6 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_5 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_4 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_3 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_2 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_1 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_0 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_5 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_5 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_5 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_4 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_4 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_4 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_3 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_3 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_3 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_2 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_2 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_2 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_1 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_1 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_1 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_0 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_0 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_0 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_93 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_92 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_91 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_90 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_89 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_88 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_87 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_86 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_85 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_84 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_83 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_82 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_81 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_80 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_79 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_78 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_77 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_76 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_75 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_74 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_73 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_72 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_71 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_70 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_69 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_68 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_67 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_66 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_65 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_64 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_63 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_62 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_61 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_60 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_59 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_58 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_57 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_56 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_55 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_54 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_53 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_52 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_51 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_50 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_49 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_48 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_47 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_46 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_45 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_44 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_43 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_42 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_41 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_40 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_39 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_38 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_37 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_36 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_35 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_34 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_33 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_32 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_31 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_30 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_29 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_28 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_27 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_26 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_25 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_24 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_23 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_22 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_21 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_20 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_19 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_18 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_17 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_16 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_15 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_14 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_13 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_12 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_11 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_10 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_9 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_8 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_7 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_6 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_5 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_4 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_3 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX4 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_2 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_1 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_0 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_30 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_29 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_28 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_27 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_26 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_25 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_24 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_23 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_22 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_21 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_20 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_19 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_18 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_17 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_16 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_15 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_14 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_13 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_12 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_11 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_10 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_9 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_8 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_7 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_6 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_5 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_4 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_3 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_2 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_1 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_0 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_30 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_131 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_130 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_129 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_128 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_29 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_127 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_126 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_125 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_124 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_28 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_123 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_122 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_121 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_120 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_27 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_119 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_118 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_117 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_116 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_26 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_115 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_114 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_113 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_112 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_25 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_111 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_110 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_109 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_108 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_24 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_107 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_106 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_105 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_104 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_23 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_103 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_102 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_101 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_100 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_22 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_99 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_98 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_97 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_96 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_21 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_95 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_94 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_93 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_92 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_20 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_91 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_90 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_89 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_88 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_19 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_87 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_86 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_85 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_84 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_18 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_83 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_82 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_81 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_80 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_17 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_79 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_78 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_77 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_76 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_16 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_75 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_74 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_73 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_72 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_15 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_71 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_70 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_69 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_68 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_14 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_67 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_66 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_65 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_64 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_13 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_63 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_62 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_61 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_60 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_12 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_59 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_58 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_57 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_56 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_11 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_55 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_54 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_53 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_52 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_10 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_51 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_50 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_49 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_48 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_9 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_47 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_46 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_45 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_44 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_8 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_43 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_42 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_41 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_40 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_7 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_39 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_38 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_37 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_36 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_6 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_35 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_34 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_33 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_32 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_5 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_31 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_30 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_29 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_28 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_4 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_27 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_26 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_25 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_24 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_3 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_23 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_22 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_21 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_20 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_2 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_19 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_18 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_17 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_16 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_1 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_15 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_14 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_13 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_12 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_0 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_11 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_10 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_9 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum) );
  evMUX2_1_8 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evlpRegister_wdt32_0 ( din, clock, reset_n, dout );
  input [31:0] din;
  output [31:0] dout;
  input clock, reset_n;


  evMS_Rstbl_FlipFlop_62 ff_0 ( .din(din[0]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[0]) );
  evMS_Rstbl_FlipFlop_61 ff_1 ( .din(din[1]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[1]) );
  evMS_Rstbl_FlipFlop_60 ff_2 ( .din(din[2]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[2]) );
  evMS_Rstbl_FlipFlop_59 ff_3 ( .din(din[3]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[3]) );
  evMS_Rstbl_FlipFlop_58 ff_4 ( .din(din[4]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[4]) );
  evMS_Rstbl_FlipFlop_57 ff_5 ( .din(din[5]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[5]) );
  evMS_Rstbl_FlipFlop_56 ff_6 ( .din(din[6]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[6]) );
  evMS_Rstbl_FlipFlop_55 ff_7 ( .din(din[7]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[7]) );
  evMS_Rstbl_FlipFlop_54 ff_8 ( .din(din[8]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[8]) );
  evMS_Rstbl_FlipFlop_53 ff_9 ( .din(din[9]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[9]) );
  evMS_Rstbl_FlipFlop_52 ff_10 ( .din(din[10]), .clock(clock), .reset_n(
        reset_n), .dout(dout[10]) );
  evMS_Rstbl_FlipFlop_51 ff_11 ( .din(din[11]), .clock(clock), .reset_n(
        reset_n), .dout(dout[11]) );
  evMS_Rstbl_FlipFlop_50 ff_12 ( .din(din[12]), .clock(clock), .reset_n(
        reset_n), .dout(dout[12]) );
  evMS_Rstbl_FlipFlop_49 ff_13 ( .din(din[13]), .clock(clock), .reset_n(
        reset_n), .dout(dout[13]) );
  evMS_Rstbl_FlipFlop_48 ff_14 ( .din(din[14]), .clock(clock), .reset_n(
        reset_n), .dout(dout[14]) );
  evMS_Rstbl_FlipFlop_47 ff_15 ( .din(din[15]), .clock(clock), .reset_n(
        reset_n), .dout(dout[15]) );
  evMS_Rstbl_FlipFlop_46 ff_16 ( .din(din[16]), .clock(clock), .reset_n(
        reset_n), .dout(dout[16]) );
  evMS_Rstbl_FlipFlop_45 ff_17 ( .din(din[17]), .clock(clock), .reset_n(
        reset_n), .dout(dout[17]) );
  evMS_Rstbl_FlipFlop_44 ff_18 ( .din(din[18]), .clock(clock), .reset_n(
        reset_n), .dout(dout[18]) );
  evMS_Rstbl_FlipFlop_43 ff_19 ( .din(din[19]), .clock(clock), .reset_n(
        reset_n), .dout(dout[19]) );
  evMS_Rstbl_FlipFlop_42 ff_20 ( .din(din[20]), .clock(clock), .reset_n(
        reset_n), .dout(dout[20]) );
  evMS_Rstbl_FlipFlop_41 ff_21 ( .din(din[21]), .clock(clock), .reset_n(
        reset_n), .dout(dout[21]) );
  evMS_Rstbl_FlipFlop_40 ff_22 ( .din(din[22]), .clock(clock), .reset_n(
        reset_n), .dout(dout[22]) );
  evMS_Rstbl_FlipFlop_39 ff_23 ( .din(din[23]), .clock(clock), .reset_n(
        reset_n), .dout(dout[23]) );
  evMS_Rstbl_FlipFlop_38 ff_24 ( .din(din[24]), .clock(clock), .reset_n(
        reset_n), .dout(dout[24]) );
  evMS_Rstbl_FlipFlop_37 ff_25 ( .din(din[25]), .clock(clock), .reset_n(
        reset_n), .dout(dout[25]) );
  evMS_Rstbl_FlipFlop_36 ff_26 ( .din(din[26]), .clock(clock), .reset_n(
        reset_n), .dout(dout[26]) );
  evMS_Rstbl_FlipFlop_35 ff_27 ( .din(din[27]), .clock(clock), .reset_n(
        reset_n), .dout(dout[27]) );
  evMS_Rstbl_FlipFlop_34 ff_28 ( .din(din[28]), .clock(clock), .reset_n(
        reset_n), .dout(dout[28]) );
  evMS_Rstbl_FlipFlop_33 ff_29 ( .din(din[29]), .clock(clock), .reset_n(
        reset_n), .dout(dout[29]) );
  evMS_Rstbl_FlipFlop_32 ff_30 ( .din(din[30]), .clock(clock), .reset_n(
        reset_n), .dout(dout[30]) );
  evMS_Rstbl_FlipFlop_31 ff_31 ( .din(din[31]), .clock(clock), .reset_n(
        reset_n), .dout(dout[31]) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_168 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X4 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_167 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_166 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_165 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_164 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_163 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_162 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_161 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_160 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_159 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_158 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_157 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_156 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_155 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_154 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_153 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_152 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_151 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_150 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_149 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_148 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_147 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_146 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_145 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_144 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_143 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_142 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_141 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_140 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_139 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_138 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_137 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  MX2XL U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_136 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_135 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_134 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_133 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_132 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_131 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_130 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_129 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_128 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_127 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_126 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_125 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_124 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_123 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_122 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_121 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_120 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_119 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_118 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_117 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_116 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_115 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_114 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_113 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_112 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_111 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_110 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_109 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_108 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_107 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_106 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_105 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_104 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_103 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_102 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_101 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_100 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_99 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_98 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_97 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_96 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_95 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_94 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_93 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_92 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_91 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_90 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_89 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_88 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_87 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_86 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_85 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_84 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_83 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_82 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_81 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_80 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_79 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_78 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_77 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_76 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_75 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_74 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_73 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_72 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_71 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_70 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_69 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_68 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_67 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_66 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_65 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_64 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_63 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_62 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_61 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_60 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_59 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_58 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_57 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_56 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_55 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_54 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_53 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_52 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_51 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_50 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_49 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_48 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_47 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_46 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_45 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_44 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_43 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_42 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_41 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_40 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_39 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_38 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_37 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_36 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_35 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_34 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_33 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_32 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_31 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_30 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_29 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_28 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_27 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_26 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_25 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_24 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_23 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_22 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_21 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_20 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_19 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_18 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_17 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_16 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_15 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_14 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_13 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_12 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_11 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_10 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_9 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_8 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_7 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_6 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_5 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_4 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_3 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_2 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_1 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_0 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X2 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evRst_Latch_cell_6 ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(reset_n), .SN(1'b1), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evPrst_Latch_cell ( din, unlock, reset_n, dout );
  input din, unlock, reset_n;
  output dout;


  TLATSRX4 dout_reg ( .G(unlock), .D(din), .RN(1'b1), .SN(reset_n), .Q(dout)
         );
endmodule


`timescale 1 ns/10 ps
module evCINV_31 ( a, a_not );
  input a;
  output a_not;


  CLKINVX1 U7 ( .A(a), .Y(a_not) );
endmodule


`timescale 1 ns/10 ps
module evLatch_cell_31 ( din, unlock, dout );
  input din, unlock;
  output dout;
  wire   n_12;
  assign n_12 = unlock;

  TLATXL dout_reg ( .G(n_12), .D(din), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evMS_Prstbl_FlipFlop ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFSX1 dout_reg ( .D(din), .CK(clock), .SN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrR_6 ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_6 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evRst_Latch_cell_6 rlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evClockGator_RngCntrP ( entr, leave, clk_in_n, rst, clk_ot );
  input entr, leave, clk_in_n, rst;
  output clk_ot;
  wire   clock_allowed, sel_lin;

  evMUX2_1_7 line_selector ( .inp1(entr), .inp2(leave), .sel(clock_allowed), 
        .mx_out(sel_lin) );
  evPrst_Latch_cell prlatch ( .din(entr), .unlock(sel_lin), .reset_n(rst), 
        .dout(clock_allowed) );
  NAND2X1 U7 ( .A(clock_allowed), .B(clk_in_n), .Y(clk_ot) );
endmodule


`timescale 1 ns/10 ps
module evMS_Rstbl_FlipFlop_94 ( din, clock, reset_n, dout );
  input din, clock, reset_n;
  output dout;


  DFFRX1 dout_reg ( .D(din), .CK(clock), .RN(reset_n), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evNMOS_31 ( src, gat, drn );
  input src, gat;
  output drn;

  tri   drn;

  TBUFX6 drn_tri ( .A(src), .OE(gat), .Y(drn) );
endmodule


`timescale 1 ns/10 ps
module evLPFA_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   a_not, a_xor_b, a_xnor_b;

  evCINV_31 inv ( .a(a), .a_not(a_not) );
  evMUX2_1_135 mx1 ( .inp1(a), .inp2(a_not), .sel(b), .mx_out(a_xor_b) );
  evMUX2_1_134 mx2 ( .inp1(a_not), .inp2(a), .sel(b), .mx_out(a_xnor_b) );
  evMUX2_1_133 mx3 ( .inp1(a_xor_b), .inp2(a_xnor_b), .sel(cin), .mx_out(sum)
         );
  evMUX2_1_132 mx4 ( .inp1(b), .inp2(cin), .sel(a_xor_b), .mx_out(cout) );
endmodule


`timescale 1 ns/10 ps
module evInpDemuxLatch_wdt32 ( din, sel, dout );
  input [31:0] sel;
  output [31:0] dout;
  input din;


  evLatch_cell_31 latch_0 ( .din(din), .unlock(sel[0]), .dout(dout[0]) );
  evLatch_cell_30 latch_1 ( .din(din), .unlock(sel[1]), .dout(dout[1]) );
  evLatch_cell_29 latch_2 ( .din(din), .unlock(sel[2]), .dout(dout[2]) );
  evLatch_cell_28 latch_3 ( .din(din), .unlock(sel[3]), .dout(dout[3]) );
  evLatch_cell_27 latch_4 ( .din(din), .unlock(sel[4]), .dout(dout[4]) );
  evLatch_cell_26 latch_5 ( .din(din), .unlock(sel[5]), .dout(dout[5]) );
  evLatch_cell_25 latch_6 ( .din(din), .unlock(sel[6]), .dout(dout[6]) );
  evLatch_cell_24 latch_7 ( .din(din), .unlock(sel[7]), .dout(dout[7]) );
  evLatch_cell_23 latch_8 ( .din(din), .unlock(sel[8]), .dout(dout[8]) );
  evLatch_cell_22 latch_9 ( .din(din), .unlock(sel[9]), .dout(dout[9]) );
  evLatch_cell_21 latch_10 ( .din(din), .unlock(sel[10]), .dout(dout[10]) );
  evLatch_cell_20 latch_11 ( .din(din), .unlock(sel[11]), .dout(dout[11]) );
  evLatch_cell_19 latch_12 ( .din(din), .unlock(sel[12]), .dout(dout[12]) );
  evLatch_cell_18 latch_13 ( .din(din), .unlock(sel[13]), .dout(dout[13]) );
  evLatch_cell_17 latch_14 ( .din(din), .unlock(sel[14]), .dout(dout[14]) );
  evLatch_cell_16 latch_15 ( .din(din), .unlock(sel[15]), .dout(dout[15]) );
  evLatch_cell_15 latch_16 ( .din(din), .unlock(sel[16]), .dout(dout[16]) );
  evLatch_cell_14 latch_17 ( .din(din), .unlock(sel[17]), .dout(dout[17]) );
  evLatch_cell_13 latch_18 ( .din(din), .unlock(sel[18]), .dout(dout[18]) );
  evLatch_cell_12 latch_19 ( .din(din), .unlock(sel[19]), .dout(dout[19]) );
  evLatch_cell_11 latch_20 ( .din(din), .unlock(sel[20]), .dout(dout[20]) );
  evLatch_cell_10 latch_21 ( .din(din), .unlock(sel[21]), .dout(dout[21]) );
  evLatch_cell_9 latch_22 ( .din(din), .unlock(sel[22]), .dout(dout[22]) );
  evLatch_cell_8 latch_23 ( .din(din), .unlock(sel[23]), .dout(dout[23]) );
  evLatch_cell_7 latch_24 ( .din(din), .unlock(sel[24]), .dout(dout[24]) );
  evLatch_cell_6 latch_25 ( .din(din), .unlock(sel[25]), .dout(dout[25]) );
  evLatch_cell_5 latch_26 ( .din(din), .unlock(sel[26]), .dout(dout[26]) );
  evLatch_cell_4 latch_27 ( .din(din), .unlock(sel[27]), .dout(dout[27]) );
  evLatch_cell_3 latch_28 ( .din(din), .unlock(sel[28]), .dout(dout[28]) );
  evLatch_cell_2 latch_29 ( .din(din), .unlock(sel[29]), .dout(dout[29]) );
  evLatch_cell_1 latch_30 ( .din(din), .unlock(sel[30]), .dout(dout[30]) );
  evLatch_cell_0 latch_31 ( .din(din), .unlock(sel[31]), .dout(dout[31]) );
endmodule


`timescale 1 ns/10 ps
module evRingCounter_GtdClk_wdt32_block_size4 ( reset_n, clock_n, dout );
  output [31:0] dout;
  input reset_n, clock_n;
  wire   \gated_clock[7] , \gated_clock[6] , \gated_clock[5] ,
         \gated_clock[4] , \gated_clock[3] , \gated_clock[2] ,
         \gated_clock[1] , \gated_clock[0] ;

  evClockGator_RngCntrP first_gator ( .entr(dout[31]), .leave(dout[4]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[0] ) );
  evClockGator_RngCntrR_6 gator_1 ( .entr(dout[3]), .leave(dout[8]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[1] ) );
  evClockGator_RngCntrR_5 gator_2 ( .entr(dout[7]), .leave(dout[12]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[2] ) );
  evClockGator_RngCntrR_4 gator_3 ( .entr(dout[11]), .leave(dout[16]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[3] ) );
  evClockGator_RngCntrR_3 gator_4 ( .entr(dout[15]), .leave(dout[20]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[4] ) );
  evClockGator_RngCntrR_2 gator_5 ( .entr(dout[19]), .leave(dout[24]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[5] ) );
  evClockGator_RngCntrR_1 gator_6 ( .entr(dout[23]), .leave(dout[28]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[6] ) );
  evClockGator_RngCntrR_0 last_gator_7 ( .entr(dout[27]), .leave(dout[0]), 
        .clk_in_n(clock_n), .rst(reset_n), .clk_ot(\gated_clock[7] ) );
  evMS_Prstbl_FlipFlop first_ff ( .din(dout[31]), .clock(\gated_clock[0] ), 
        .reset_n(reset_n), .dout(dout[0]) );
  evMS_Rstbl_FlipFlop_30 ff_1 ( .din(dout[0]), .clock(\gated_clock[0] ), 
        .reset_n(reset_n), .dout(dout[1]) );
  evMS_Rstbl_FlipFlop_29 ff_2 ( .din(dout[1]), .clock(\gated_clock[0] ), 
        .reset_n(reset_n), .dout(dout[2]) );
  evMS_Rstbl_FlipFlop_28 ff_3 ( .din(dout[2]), .clock(\gated_clock[0] ), 
        .reset_n(reset_n), .dout(dout[3]) );
  evMS_Rstbl_FlipFlop_27 ff_4 ( .din(dout[3]), .clock(\gated_clock[1] ), 
        .reset_n(reset_n), .dout(dout[4]) );
  evMS_Rstbl_FlipFlop_26 ff_5 ( .din(dout[4]), .clock(\gated_clock[1] ), 
        .reset_n(reset_n), .dout(dout[5]) );
  evMS_Rstbl_FlipFlop_25 ff_6 ( .din(dout[5]), .clock(\gated_clock[1] ), 
        .reset_n(reset_n), .dout(dout[6]) );
  evMS_Rstbl_FlipFlop_24 ff_7 ( .din(dout[6]), .clock(\gated_clock[1] ), 
        .reset_n(reset_n), .dout(dout[7]) );
  evMS_Rstbl_FlipFlop_23 ff_8 ( .din(dout[7]), .clock(\gated_clock[2] ), 
        .reset_n(reset_n), .dout(dout[8]) );
  evMS_Rstbl_FlipFlop_22 ff_9 ( .din(dout[8]), .clock(\gated_clock[2] ), 
        .reset_n(reset_n), .dout(dout[9]) );
  evMS_Rstbl_FlipFlop_21 ff_10 ( .din(dout[9]), .clock(\gated_clock[2] ), 
        .reset_n(reset_n), .dout(dout[10]) );
  evMS_Rstbl_FlipFlop_20 ff_11 ( .din(dout[10]), .clock(\gated_clock[2] ), 
        .reset_n(reset_n), .dout(dout[11]) );
  evMS_Rstbl_FlipFlop_19 ff_12 ( .din(dout[11]), .clock(\gated_clock[3] ), 
        .reset_n(reset_n), .dout(dout[12]) );
  evMS_Rstbl_FlipFlop_18 ff_13 ( .din(dout[12]), .clock(\gated_clock[3] ), 
        .reset_n(reset_n), .dout(dout[13]) );
  evMS_Rstbl_FlipFlop_17 ff_14 ( .din(dout[13]), .clock(\gated_clock[3] ), 
        .reset_n(reset_n), .dout(dout[14]) );
  evMS_Rstbl_FlipFlop_16 ff_15 ( .din(dout[14]), .clock(\gated_clock[3] ), 
        .reset_n(reset_n), .dout(dout[15]) );
  evMS_Rstbl_FlipFlop_15 ff_16 ( .din(dout[15]), .clock(\gated_clock[4] ), 
        .reset_n(reset_n), .dout(dout[16]) );
  evMS_Rstbl_FlipFlop_14 ff_17 ( .din(dout[16]), .clock(\gated_clock[4] ), 
        .reset_n(reset_n), .dout(dout[17]) );
  evMS_Rstbl_FlipFlop_13 ff_18 ( .din(dout[17]), .clock(\gated_clock[4] ), 
        .reset_n(reset_n), .dout(dout[18]) );
  evMS_Rstbl_FlipFlop_12 ff_19 ( .din(dout[18]), .clock(\gated_clock[4] ), 
        .reset_n(reset_n), .dout(dout[19]) );
  evMS_Rstbl_FlipFlop_11 ff_20 ( .din(dout[19]), .clock(\gated_clock[5] ), 
        .reset_n(reset_n), .dout(dout[20]) );
  evMS_Rstbl_FlipFlop_10 ff_21 ( .din(dout[20]), .clock(\gated_clock[5] ), 
        .reset_n(reset_n), .dout(dout[21]) );
  evMS_Rstbl_FlipFlop_9 ff_22 ( .din(dout[21]), .clock(\gated_clock[5] ), 
        .reset_n(reset_n), .dout(dout[22]) );
  evMS_Rstbl_FlipFlop_8 ff_23 ( .din(dout[22]), .clock(\gated_clock[5] ), 
        .reset_n(reset_n), .dout(dout[23]) );
  evMS_Rstbl_FlipFlop_7 ff_24 ( .din(dout[23]), .clock(\gated_clock[6] ), 
        .reset_n(reset_n), .dout(dout[24]) );
  evMS_Rstbl_FlipFlop_6 ff_25 ( .din(dout[24]), .clock(\gated_clock[6] ), 
        .reset_n(reset_n), .dout(dout[25]) );
  evMS_Rstbl_FlipFlop_5 ff_26 ( .din(dout[25]), .clock(\gated_clock[6] ), 
        .reset_n(reset_n), .dout(dout[26]) );
  evMS_Rstbl_FlipFlop_4 ff_27 ( .din(dout[26]), .clock(\gated_clock[6] ), 
        .reset_n(reset_n), .dout(dout[27]) );
  evMS_Rstbl_FlipFlop_3 ff_28 ( .din(dout[27]), .clock(\gated_clock[7] ), 
        .reset_n(reset_n), .dout(dout[28]) );
  evMS_Rstbl_FlipFlop_2 ff_29 ( .din(dout[28]), .clock(\gated_clock[7] ), 
        .reset_n(reset_n), .dout(dout[29]) );
  evMS_Rstbl_FlipFlop_1 ff_30 ( .din(dout[29]), .clock(\gated_clock[7] ), 
        .reset_n(reset_n), .dout(dout[30]) );
  evMS_Rstbl_FlipFlop_0 ff_31 ( .din(dout[30]), .clock(\gated_clock[7] ), 
        .reset_n(reset_n), .dout(dout[31]) );
endmodule


`timescale 1 ns/10 ps
module evlpMux2_1_wdt33 ( inp1, inp2, sel, mx_out );
  input [32:0] inp1;
  input [32:0] inp2;
  output [32:0] mx_out;
  input sel;


  evMUX2_1_168 mux_0 ( .inp1(inp1[0]), .inp2(inp2[0]), .sel(sel), .mx_out(
        mx_out[0]) );
  evMUX2_1_167 mux_1 ( .inp1(inp1[1]), .inp2(inp2[1]), .sel(sel), .mx_out(
        mx_out[1]) );
  evMUX2_1_166 mux_2 ( .inp1(inp1[2]), .inp2(inp2[2]), .sel(sel), .mx_out(
        mx_out[2]) );
  evMUX2_1_165 mux_3 ( .inp1(inp1[3]), .inp2(inp2[3]), .sel(sel), .mx_out(
        mx_out[3]) );
  evMUX2_1_164 mux_4 ( .inp1(inp1[4]), .inp2(inp2[4]), .sel(sel), .mx_out(
        mx_out[4]) );
  evMUX2_1_163 mux_5 ( .inp1(inp1[5]), .inp2(inp2[5]), .sel(sel), .mx_out(
        mx_out[5]) );
  evMUX2_1_162 mux_6 ( .inp1(inp1[6]), .inp2(inp2[6]), .sel(sel), .mx_out(
        mx_out[6]) );
  evMUX2_1_161 mux_7 ( .inp1(inp1[7]), .inp2(inp2[7]), .sel(sel), .mx_out(
        mx_out[7]) );
  evMUX2_1_160 mux_8 ( .inp1(inp1[8]), .inp2(inp2[8]), .sel(sel), .mx_out(
        mx_out[8]) );
  evMUX2_1_159 mux_9 ( .inp1(inp1[9]), .inp2(inp2[9]), .sel(sel), .mx_out(
        mx_out[9]) );
  evMUX2_1_158 mux_10 ( .inp1(inp1[10]), .inp2(inp2[10]), .sel(sel), .mx_out(
        mx_out[10]) );
  evMUX2_1_157 mux_11 ( .inp1(inp1[11]), .inp2(inp2[11]), .sel(sel), .mx_out(
        mx_out[11]) );
  evMUX2_1_156 mux_12 ( .inp1(inp1[12]), .inp2(inp2[12]), .sel(sel), .mx_out(
        mx_out[12]) );
  evMUX2_1_155 mux_13 ( .inp1(inp1[13]), .inp2(inp2[13]), .sel(sel), .mx_out(
        mx_out[13]) );
  evMUX2_1_154 mux_14 ( .inp1(inp1[14]), .inp2(inp2[14]), .sel(sel), .mx_out(
        mx_out[14]) );
  evMUX2_1_153 mux_15 ( .inp1(inp1[15]), .inp2(inp2[15]), .sel(sel), .mx_out(
        mx_out[15]) );
  evMUX2_1_152 mux_16 ( .inp1(inp1[16]), .inp2(inp2[16]), .sel(sel), .mx_out(
        mx_out[16]) );
  evMUX2_1_151 mux_17 ( .inp1(inp1[17]), .inp2(inp2[17]), .sel(sel), .mx_out(
        mx_out[17]) );
  evMUX2_1_150 mux_18 ( .inp1(inp1[18]), .inp2(inp2[18]), .sel(sel), .mx_out(
        mx_out[18]) );
  evMUX2_1_149 mux_19 ( .inp1(inp1[19]), .inp2(inp2[19]), .sel(sel), .mx_out(
        mx_out[19]) );
  evMUX2_1_148 mux_20 ( .inp1(inp1[20]), .inp2(inp2[20]), .sel(sel), .mx_out(
        mx_out[20]) );
  evMUX2_1_147 mux_21 ( .inp1(inp1[21]), .inp2(inp2[21]), .sel(sel), .mx_out(
        mx_out[21]) );
  evMUX2_1_146 mux_22 ( .inp1(inp1[22]), .inp2(inp2[22]), .sel(sel), .mx_out(
        mx_out[22]) );
  evMUX2_1_145 mux_23 ( .inp1(inp1[23]), .inp2(inp2[23]), .sel(sel), .mx_out(
        mx_out[23]) );
  evMUX2_1_144 mux_24 ( .inp1(inp1[24]), .inp2(inp2[24]), .sel(sel), .mx_out(
        mx_out[24]) );
  evMUX2_1_143 mux_25 ( .inp1(inp1[25]), .inp2(inp2[25]), .sel(sel), .mx_out(
        mx_out[25]) );
  evMUX2_1_142 mux_26 ( .inp1(inp1[26]), .inp2(inp2[26]), .sel(sel), .mx_out(
        mx_out[26]) );
  evMUX2_1_141 mux_27 ( .inp1(inp1[27]), .inp2(inp2[27]), .sel(sel), .mx_out(
        mx_out[27]) );
  evMUX2_1_140 mux_28 ( .inp1(inp1[28]), .inp2(inp2[28]), .sel(sel), .mx_out(
        mx_out[28]) );
  evMUX2_1_139 mux_29 ( .inp1(inp1[29]), .inp2(inp2[29]), .sel(sel), .mx_out(
        mx_out[29]) );
  evMUX2_1_138 mux_30 ( .inp1(inp1[30]), .inp2(inp2[30]), .sel(sel), .mx_out(
        mx_out[30]) );
  evMUX2_1_137 mux_31 ( .inp1(inp1[31]), .inp2(inp2[31]), .sel(sel), .mx_out(
        mx_out[31]) );
  evMUX2_1_136 mux_32 ( .inp1(inp1[32]), .inp2(inp2[32]), .sel(sel), .mx_out(
        mx_out[32]) );
endmodule


`timescale 1 ns/10 ps
module evlpRegister_wdt32_1 ( din, clock, reset_n, dout );
  input [31:0] din;
  output [31:0] dout;
  input clock, reset_n;


  evMS_Rstbl_FlipFlop_94 ff_0 ( .din(din[0]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[0]) );
  evMS_Rstbl_FlipFlop_93 ff_1 ( .din(din[1]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[1]) );
  evMS_Rstbl_FlipFlop_92 ff_2 ( .din(din[2]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[2]) );
  evMS_Rstbl_FlipFlop_91 ff_3 ( .din(din[3]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[3]) );
  evMS_Rstbl_FlipFlop_90 ff_4 ( .din(din[4]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[4]) );
  evMS_Rstbl_FlipFlop_89 ff_5 ( .din(din[5]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[5]) );
  evMS_Rstbl_FlipFlop_88 ff_6 ( .din(din[6]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[6]) );
  evMS_Rstbl_FlipFlop_87 ff_7 ( .din(din[7]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[7]) );
  evMS_Rstbl_FlipFlop_86 ff_8 ( .din(din[8]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[8]) );
  evMS_Rstbl_FlipFlop_85 ff_9 ( .din(din[9]), .clock(clock), .reset_n(reset_n), 
        .dout(dout[9]) );
  evMS_Rstbl_FlipFlop_84 ff_10 ( .din(din[10]), .clock(clock), .reset_n(
        reset_n), .dout(dout[10]) );
  evMS_Rstbl_FlipFlop_83 ff_11 ( .din(din[11]), .clock(clock), .reset_n(
        reset_n), .dout(dout[11]) );
  evMS_Rstbl_FlipFlop_82 ff_12 ( .din(din[12]), .clock(clock), .reset_n(
        reset_n), .dout(dout[12]) );
  evMS_Rstbl_FlipFlop_81 ff_13 ( .din(din[13]), .clock(clock), .reset_n(
        reset_n), .dout(dout[13]) );
  evMS_Rstbl_FlipFlop_80 ff_14 ( .din(din[14]), .clock(clock), .reset_n(
        reset_n), .dout(dout[14]) );
  evMS_Rstbl_FlipFlop_79 ff_15 ( .din(din[15]), .clock(clock), .reset_n(
        reset_n), .dout(dout[15]) );
  evMS_Rstbl_FlipFlop_78 ff_16 ( .din(din[16]), .clock(clock), .reset_n(
        reset_n), .dout(dout[16]) );
  evMS_Rstbl_FlipFlop_77 ff_17 ( .din(din[17]), .clock(clock), .reset_n(
        reset_n), .dout(dout[17]) );
  evMS_Rstbl_FlipFlop_76 ff_18 ( .din(din[18]), .clock(clock), .reset_n(
        reset_n), .dout(dout[18]) );
  evMS_Rstbl_FlipFlop_75 ff_19 ( .din(din[19]), .clock(clock), .reset_n(
        reset_n), .dout(dout[19]) );
  evMS_Rstbl_FlipFlop_74 ff_20 ( .din(din[20]), .clock(clock), .reset_n(
        reset_n), .dout(dout[20]) );
  evMS_Rstbl_FlipFlop_73 ff_21 ( .din(din[21]), .clock(clock), .reset_n(
        reset_n), .dout(dout[21]) );
  evMS_Rstbl_FlipFlop_72 ff_22 ( .din(din[22]), .clock(clock), .reset_n(
        reset_n), .dout(dout[22]) );
  evMS_Rstbl_FlipFlop_71 ff_23 ( .din(din[23]), .clock(clock), .reset_n(
        reset_n), .dout(dout[23]) );
  evMS_Rstbl_FlipFlop_70 ff_24 ( .din(din[24]), .clock(clock), .reset_n(
        reset_n), .dout(dout[24]) );
  evMS_Rstbl_FlipFlop_69 ff_25 ( .din(din[25]), .clock(clock), .reset_n(
        reset_n), .dout(dout[25]) );
  evMS_Rstbl_FlipFlop_68 ff_26 ( .din(din[26]), .clock(clock), .reset_n(
        reset_n), .dout(dout[26]) );
  evMS_Rstbl_FlipFlop_67 ff_27 ( .din(din[27]), .clock(clock), .reset_n(
        reset_n), .dout(dout[27]) );
  evMS_Rstbl_FlipFlop_66 ff_28 ( .din(din[28]), .clock(clock), .reset_n(
        reset_n), .dout(dout[28]) );
  evMS_Rstbl_FlipFlop_65 ff_29 ( .din(din[29]), .clock(clock), .reset_n(
        reset_n), .dout(dout[29]) );
  evMS_Rstbl_FlipFlop_64 ff_30 ( .din(din[30]), .clock(clock), .reset_n(
        reset_n), .dout(dout[30]) );
  evMS_Rstbl_FlipFlop_63 ff_31 ( .din(din[31]), .clock(clock), .reset_n(
        reset_n), .dout(dout[31]) );
endmodule


`timescale 1 ns/10 ps
module evNonEncodedMux_wdt32 ( din, sel, dout );
  input [31:0] din;
  input [31:0] sel;
  output dout;

  tri   dout;

  evNMOS_31 nms_0 ( .src(din[0]), .gat(sel[0]), .drn(dout) );
  evNMOS_30 nms_1 ( .src(din[1]), .gat(sel[1]), .drn(dout) );
  evNMOS_29 nms_2 ( .src(din[2]), .gat(sel[2]), .drn(dout) );
  evNMOS_28 nms_3 ( .src(din[3]), .gat(sel[3]), .drn(dout) );
  evNMOS_27 nms_4 ( .src(din[4]), .gat(sel[4]), .drn(dout) );
  evNMOS_26 nms_5 ( .src(din[5]), .gat(sel[5]), .drn(dout) );
  evNMOS_25 nms_6 ( .src(din[6]), .gat(sel[6]), .drn(dout) );
  evNMOS_24 nms_7 ( .src(din[7]), .gat(sel[7]), .drn(dout) );
  evNMOS_23 nms_8 ( .src(din[8]), .gat(sel[8]), .drn(dout) );
  evNMOS_22 nms_9 ( .src(din[9]), .gat(sel[9]), .drn(dout) );
  evNMOS_21 nms_10 ( .src(din[10]), .gat(sel[10]), .drn(dout) );
  evNMOS_20 nms_11 ( .src(din[11]), .gat(sel[11]), .drn(dout) );
  evNMOS_19 nms_12 ( .src(din[12]), .gat(sel[12]), .drn(dout) );
  evNMOS_18 nms_13 ( .src(din[13]), .gat(sel[13]), .drn(dout) );
  evNMOS_17 nms_14 ( .src(din[14]), .gat(sel[14]), .drn(dout) );
  evNMOS_16 nms_15 ( .src(din[15]), .gat(sel[15]), .drn(dout) );
  evNMOS_15 nms_16 ( .src(din[16]), .gat(sel[16]), .drn(dout) );
  evNMOS_14 nms_17 ( .src(din[17]), .gat(sel[17]), .drn(dout) );
  evNMOS_13 nms_18 ( .src(din[18]), .gat(sel[18]), .drn(dout) );
  evNMOS_12 nms_19 ( .src(din[19]), .gat(sel[19]), .drn(dout) );
  evNMOS_11 nms_20 ( .src(din[20]), .gat(sel[20]), .drn(dout) );
  evNMOS_10 nms_21 ( .src(din[21]), .gat(sel[21]), .drn(dout) );
  evNMOS_9 nms_22 ( .src(din[22]), .gat(sel[22]), .drn(dout) );
  evNMOS_8 nms_23 ( .src(din[23]), .gat(sel[23]), .drn(dout) );
  evNMOS_7 nms_24 ( .src(din[24]), .gat(sel[24]), .drn(dout) );
  evNMOS_6 nms_25 ( .src(din[25]), .gat(sel[25]), .drn(dout) );
  evNMOS_5 nms_26 ( .src(din[26]), .gat(sel[26]), .drn(dout) );
  evNMOS_4 nms_27 ( .src(din[27]), .gat(sel[27]), .drn(dout) );
  evNMOS_3 nms_28 ( .src(din[28]), .gat(sel[28]), .drn(dout) );
  evNMOS_2 nms_29 ( .src(din[29]), .gat(sel[29]), .drn(dout) );
  evNMOS_1 nms_30 ( .src(din[30]), .gat(sel[30]), .drn(dout) );
  evNMOS_0 nms_31 ( .src(din[31]), .gat(sel[31]), .drn(dout) );
endmodule


`timescale 1 ns/10 ps
module evlpRCAdder_wdt32 ( a, b, cin, sum, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout;
  wire   \imsg[31] , \imsg[30] , \imsg[29] , \imsg[28] , \imsg[27] ,
         \imsg[26] , \imsg[25] , \imsg[24] , \imsg[23] , \imsg[22] ,
         \imsg[21] , \imsg[20] , \imsg[19] , \imsg[18] , \imsg[17] ,
         \imsg[16] , \imsg[15] , \imsg[14] , \imsg[13] , \imsg[12] ,
         \imsg[11] , \imsg[10] , \imsg[9] , \imsg[8] , \imsg[7] , \imsg[6] ,
         \imsg[5] , \imsg[4] , \imsg[3] , \imsg[2] , \imsg[1] ;

  evLPFA_31 adder_0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        \imsg[1] ) );
  evLPFA_30 adder_1 ( .a(a[1]), .b(b[1]), .cin(\imsg[1] ), .sum(sum[1]), 
        .cout(\imsg[2] ) );
  evLPFA_29 adder_2 ( .a(a[2]), .b(b[2]), .cin(\imsg[2] ), .sum(sum[2]), 
        .cout(\imsg[3] ) );
  evLPFA_28 adder_3 ( .a(a[3]), .b(b[3]), .cin(\imsg[3] ), .sum(sum[3]), 
        .cout(\imsg[4] ) );
  evLPFA_27 adder_4 ( .a(a[4]), .b(b[4]), .cin(\imsg[4] ), .sum(sum[4]), 
        .cout(\imsg[5] ) );
  evLPFA_26 adder_5 ( .a(a[5]), .b(b[5]), .cin(\imsg[5] ), .sum(sum[5]), 
        .cout(\imsg[6] ) );
  evLPFA_25 adder_6 ( .a(a[6]), .b(b[6]), .cin(\imsg[6] ), .sum(sum[6]), 
        .cout(\imsg[7] ) );
  evLPFA_24 adder_7 ( .a(a[7]), .b(b[7]), .cin(\imsg[7] ), .sum(sum[7]), 
        .cout(\imsg[8] ) );
  evLPFA_23 adder_8 ( .a(a[8]), .b(b[8]), .cin(\imsg[8] ), .sum(sum[8]), 
        .cout(\imsg[9] ) );
  evLPFA_22 adder_9 ( .a(a[9]), .b(b[9]), .cin(\imsg[9] ), .sum(sum[9]), 
        .cout(\imsg[10] ) );
  evLPFA_21 adder_10 ( .a(a[10]), .b(b[10]), .cin(\imsg[10] ), .sum(sum[10]), 
        .cout(\imsg[11] ) );
  evLPFA_20 adder_11 ( .a(a[11]), .b(b[11]), .cin(\imsg[11] ), .sum(sum[11]), 
        .cout(\imsg[12] ) );
  evLPFA_19 adder_12 ( .a(a[12]), .b(b[12]), .cin(\imsg[12] ), .sum(sum[12]), 
        .cout(\imsg[13] ) );
  evLPFA_18 adder_13 ( .a(a[13]), .b(b[13]), .cin(\imsg[13] ), .sum(sum[13]), 
        .cout(\imsg[14] ) );
  evLPFA_17 adder_14 ( .a(a[14]), .b(b[14]), .cin(\imsg[14] ), .sum(sum[14]), 
        .cout(\imsg[15] ) );
  evLPFA_16 adder_15 ( .a(a[15]), .b(b[15]), .cin(\imsg[15] ), .sum(sum[15]), 
        .cout(\imsg[16] ) );
  evLPFA_15 adder_16 ( .a(a[16]), .b(b[16]), .cin(\imsg[16] ), .sum(sum[16]), 
        .cout(\imsg[17] ) );
  evLPFA_14 adder_17 ( .a(a[17]), .b(b[17]), .cin(\imsg[17] ), .sum(sum[17]), 
        .cout(\imsg[18] ) );
  evLPFA_13 adder_18 ( .a(a[18]), .b(b[18]), .cin(\imsg[18] ), .sum(sum[18]), 
        .cout(\imsg[19] ) );
  evLPFA_12 adder_19 ( .a(a[19]), .b(b[19]), .cin(\imsg[19] ), .sum(sum[19]), 
        .cout(\imsg[20] ) );
  evLPFA_11 adder_20 ( .a(a[20]), .b(b[20]), .cin(\imsg[20] ), .sum(sum[20]), 
        .cout(\imsg[21] ) );
  evLPFA_10 adder_21 ( .a(a[21]), .b(b[21]), .cin(\imsg[21] ), .sum(sum[21]), 
        .cout(\imsg[22] ) );
  evLPFA_9 adder_22 ( .a(a[22]), .b(b[22]), .cin(\imsg[22] ), .sum(sum[22]), 
        .cout(\imsg[23] ) );
  evLPFA_8 adder_23 ( .a(a[23]), .b(b[23]), .cin(\imsg[23] ), .sum(sum[23]), 
        .cout(\imsg[24] ) );
  evLPFA_7 adder_24 ( .a(a[24]), .b(b[24]), .cin(\imsg[24] ), .sum(sum[24]), 
        .cout(\imsg[25] ) );
  evLPFA_6 adder_25 ( .a(a[25]), .b(b[25]), .cin(\imsg[25] ), .sum(sum[25]), 
        .cout(\imsg[26] ) );
  evLPFA_5 adder_26 ( .a(a[26]), .b(b[26]), .cin(\imsg[26] ), .sum(sum[26]), 
        .cout(\imsg[27] ) );
  evLPFA_4 adder_27 ( .a(a[27]), .b(b[27]), .cin(\imsg[27] ), .sum(sum[27]), 
        .cout(\imsg[28] ) );
  evLPFA_3 adder_28 ( .a(a[28]), .b(b[28]), .cin(\imsg[28] ), .sum(sum[28]), 
        .cout(\imsg[29] ) );
  evLPFA_2 adder_29 ( .a(a[29]), .b(b[29]), .cin(\imsg[29] ), .sum(sum[29]), 
        .cout(\imsg[30] ) );
  evLPFA_1 adder_30 ( .a(a[30]), .b(b[30]), .cin(\imsg[30] ), .sum(sum[30]), 
        .cout(\imsg[31] ) );
  evLPFA_0 adder_31 ( .a(a[31]), .b(b[31]), .cin(\imsg[31] ), .sum(sum[31]), 
        .cout(cout) );
endmodule


`timescale 1 ns/10 ps
module evMUX2_1_169 ( inp1, inp2, sel, mx_out );
  input inp1, inp2, sel;
  output mx_out;


  CLKMX2X4 U10 ( .A(inp1), .B(inp2), .S0(sel), .Y(mx_out) );
endmodule


`timescale 1 ns/10 ps
module evMS_FlipFlop ( din, clock, dout );
  input din, clock;
  output dout;

  tri   din;

  DFFQX1 dout_reg ( .D(din), .CK(clock), .Q(dout) );
endmodule


`timescale 1 ns/10 ps
module evlpMultiplier ( a, b, rst, clk, clk_n, res );
  input [31:0] a;
  input [31:0] b;
  output [63:0] res;
  input rst, clk, clk_n;
  wire   bypreg_clk, fedreg_clk, cout, \this_cycle_result[0] , hot_B_bit,
         data_source_selector;
  wire   [31:0] adder_out;
  wire   [31:0] bypassed_operand;
  wire   [31:0] hot_bit_selector;
  wire   [31:0] adder_2nd_inp;
  tri   next_hot_B_bit;

  evMS_FlipFlop hot_B_bit_ff ( .din(next_hot_B_bit), .clock(clk), .dout(
        hot_B_bit) );
  evMUX2_1_169 src_sel_mux ( .inp1(hot_B_bit), .inp2(b[0]), .sel(
        hot_bit_selector[0]), .mx_out(data_source_selector) );
  evlpRCAdder_wdt32 adder ( .a(a), .b(adder_2nd_inp), .cin(1'b0), .sum(
        adder_out), .cout(cout) );
  evNonEncodedMux_wdt32 nxt_hot_bit_mux ( .din({1'b0, b[31:1]}), .sel(
        hot_bit_selector), .dout(next_hot_B_bit) );
  evlpRegister_wdt32_1 bypass_reg ( .din(res[63:32]), .clock(bypreg_clk), 
        .reset_n(rst), .dout(bypassed_operand) );
  evlpRegister_wdt32_0 feeder_reg ( .din(res[63:32]), .clock(fedreg_clk), 
        .reset_n(rst), .dout(adder_2nd_inp) );
  evlpMux2_1_wdt33 mux ( .inp1({1'b0, bypassed_operand}), .inp2({cout, 
        adder_out}), .sel(data_source_selector), .mx_out({res[63:32], 
        \this_cycle_result[0] }) );
  evRingCounter_GtdClk_wdt32_block_size4 counter ( .reset_n(rst), .clock_n(
        clk_n), .dout(hot_bit_selector) );
  evInpDemuxLatch_wdt32 low_res_latch ( .din(\this_cycle_result[0] ), .sel(
        hot_bit_selector), .dout(res[31:0]) );
  NAND2X4 U8 ( .A(next_hot_B_bit), .B(clk_n), .Y(fedreg_clk) );
  NOR2X4 U9 ( .A(next_hot_B_bit), .B(clk_n), .Y(bypreg_clk) );
endmodule

